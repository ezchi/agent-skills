module {{module_name}} #(
  parameter integer P_WIDTH = {{width}}
)(
  input  logic iClk,
  input  logic iRst,
  input  logic [P_WIDTH-1:0] iData,
  output logic [P_WIDTH-1:0] oData
);

  // TODO: Insert combinational logic here
  // TODO: Insert sequential logic here

endmodule
