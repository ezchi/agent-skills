module {{module_name}} #(
  parameter integer P_WIDTH = {{width}}
)(
  input  logic i_clk_core,
  input  logic i_rst_core,
  input  logic [P_WIDTH-1:0] i_din,
  output logic [P_WIDTH-1:0] o_dout
);

  // TODO: Insert combinational logic here
  // TODO: Insert sequential logic here

endmodule
